
always @(state ,x)
	begin
		case(state)
			A:
				begin
					if(x==0)
						next_state<=E;
					else
						next_state<=D;
			B:
				begin
					if(x==0)
						next_state<=F;
					else
						next_state<=D;
			C:
				begin
					if(x==0)
						next_state<=E;
					else
						next_state<=B;
			D:
				begin
					if(x==0)
						next_state<=F;
					else
						next_state<=B;
			E:
				begin
					if(x==0)
						next_state<=C;
					else
						next_state<=F;
			F:
				begin
					if(x==0)
						next_state<=B;
					else
						next_state<=C;
		endcase
	end
